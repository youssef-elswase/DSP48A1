module DSP48A1 #(parameter A0REG = 0 , A1REG = 1,B0REG = 0 , B1REG = 1,
    CREG = 1 ,DREG = 1,MREG = 1 ,PREG = 1,CARRYINREG = 1 ,CARRYOUTREG = 1,OPMODEREG = 1,
    CARRYINSEL = "OPMODE5" , // OPMODE5 OR CARRYIN
    B_INPUT = "DIRECT" , // DIRECT OR CASCADE
    RSTTYPR = "SYNC"  //ASYNC OR SYNC
    ) (A,B,C,D,BCIN,CARRYIN,M,P,CARRYOUT,CARRYOUTF,CLK,OPMODE,
    CEA,CEB,CEC,CECARRYIN,CED,CEM,CEOPMODE,CEP,
    RSTA,RSTB,RSTC,RSTCARRYIN,RSTD,RSTM,RSTOPMODE,RSTP,
    BCOUT,PCIN,PCOUT);

    input [17:0] A,B,D,BCIN;
    input [47:0] C,PCIN;
    input [7:0] OPMODE;
    input CARRYIN,CEA,CEB,CEC,CECARRYIN,CED,CEM,CEOPMODE,CEP,RSTA,RSTB,RSTC,RSTCARRYIN,RSTD,RSTM,RSTOPMODE,RSTP,CLK;
    output [35:0] M;
    output [47:0] P;
    output [47:0] PCOUT;
    output [17:0] BCOUT;
    output CARRYOUT;
    output CARRYOUTF;
    wire [17:0] B_IN,MDO,MB0O,MB1O,MA0O,MA1O,PREO,MADDO,AOUT;
    wire [47:0] MULO,MCO,XOUT,ZOUT,POSTO,DAB;
    wire CY0O,CY0IN,CY1O,CY1IN;
    wire [7:0] OPMODEO;
    wire [47:0] MOUT;



    REG_MUL #(RSTTYPR,1) op0 (OPMODEREG,OPMODE[0],OPMODEO[0],CLK,RSTOPMODE,CEOPMODE);
    REG_MUL #(RSTTYPR,1) op1 (OPMODEREG,OPMODE[1],OPMODEO[1],CLK,RSTOPMODE,CEOPMODE);
    REG_MUL #(RSTTYPR,1) op2 (OPMODEREG,OPMODE[2],OPMODEO[2],CLK,RSTOPMODE,CEOPMODE);
    REG_MUL #(RSTTYPR,1) op3 (OPMODEREG,OPMODE[3],OPMODEO[3],CLK,RSTOPMODE,CEOPMODE);
    REG_MUL #(RSTTYPR,1) op4 (OPMODEREG,OPMODE[4],OPMODEO[4],CLK,RSTOPMODE,CEOPMODE);
    REG_MUL #(RSTTYPR,1) op5 (OPMODEREG,OPMODE[5],OPMODEO[5],CLK,RSTOPMODE,CEOPMODE);
    REG_MUL #(RSTTYPR,1) op6 (OPMODEREG,OPMODE[6],OPMODEO[6],CLK,RSTOPMODE,CEOPMODE);
    REG_MUL #(RSTTYPR,1) op7 (OPMODEREG,OPMODE[7],OPMODEO[7],CLK,RSTOPMODE,CEOPMODE);
    assign B_IN = (B_INPUT == "DIRECT") ? B     : 
                  (B_INPUT == "CASCADE") ? BCIN : 0 ;
    REG_MUL #(RSTTYPR,18) D_r (DREG,D,MDO,CLK,RSTD,CED);
    REG_MUL #(RSTTYPR,18) B0 (B0REG,B_IN,MB0O,CLK,RSTB,CEB);
    REG_MUL #(RSTTYPR,18) A0 (A0REG,A,MA0O,CLK,RSTA,CEA);
    REG_MUL #(RSTTYPR,48) C_r (CREG,C,MCO,CLK,RSTC,CEC);
    ADD_SUB_PRE #(18) ADD_SUB1 (MDO,MB0O,PREO,OPMODEO[6]);
    assign MADDO = (OPMODEO[4]) ? PREO : MB0O ;
    REG_MUL #(RSTTYPR,18) B1 (B1REG,MADDO,BCOUT,CLK,RSTB,CEB);
    REG_MUL #(RSTTYPR,18) A1 (A1REG,MA0O,AOUT,CLK,RSTA,CEA);
    MUL #(18) MULT (BCOUT,AOUT,MULO);
    assign M = MOUT[36:0];
    REG_MUL #(RSTTYPR,48) M_r (MREG,MULO,MOUT,CLK,RSTM,CEM);
    assign DAB = {D[11:0],AOUT,BCOUT};
    assign XOUT = (OPMODEO[1:0] == 0) ? 0 :
                  (OPMODEO[1:0] == 1) ? {12'h000,M} :
                  (OPMODEO[1:0] == 2) ? P : 
                  (OPMODEO[1:0] == 3) ? DAB : 0 ;
    assign ZOUT = (OPMODEO[3:2] == 0) ? 0 :
                  (OPMODEO[3:2] == 1) ? PCIN :
                  (OPMODEO[3:2] == 2) ? P : 
                  (OPMODEO[3:2] == 3) ? MCO : 0 ;
    assign CY1IN = (CARRYINSEL == "OPMODE5") ? OPMODEO[5] : 
                   (CARRYINSEL == "CARRYIN") ? CARRYIN    : 0 ; 
    REG_MUL #(RSTTYPR,1) CY1 (CARRYINREG,CY1IN,CY1O,CLK,RSTCARRYIN,CECARRYIN);
    ADD_SUB_POST #(48) ADD_SUB2 (XOUT,ZOUT,POSTO,OPMODEO[7],CY1IN,CY0IN);
    REG_MUL #(RSTTYPR,1) CY0 (CARRYOUTREG,CY0IN,CARRYOUT,CLK,RSTCARRYIN,CECARRYIN);
    REG_MUL #(RSTTYPR,48) P_r (PREG,POSTO,P,CLK,RSTP,CEP);
    assign PCOUT = P;
    assign CARRYOUTF = CARRYOUT;

 endmodule